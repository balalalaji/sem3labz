`timescale 1ns/1ns
`include "q1.v"
module q1_tb();
reg a,b,x,y,s0,s1;
wire f;
q1 qu(s);