`timescale 1ns/1ns
`include "qtwo.v"
module qtwo_tb();
reg a,b,c,d;
wire f,g;
qtwo qu2(a,b,c,d,f,g);
initial
begin
$dumpfile("qtwo_tb.vcd");
$dumpvars(0, qtwo_tb);
	a=1'b0; b=1'b0; c=1'b0; d=1'b0; #20;
	a=1'b0; b=1'b0; c=1'b0; d=1'b1; #20;
	a=1'b0; b=1'b0; c=1'b1; d=1'b0; #20;
	a=1'b0; b=1'b0; c=1'b1; d=1'b1; #20;
	a=1'b0; b=1'b1; c=1'b0; d=1'b0; #20;
	a=1'b0; b=1'b1; c=1'b0; d=1'b1; #20;
	a=1'b0; b=1'b1; c=1'b1; d=1'b0; #20;	
	a=1'b0; b=1'b1; c=1'b1; d=1'b1; #20;
	a=1'b0; b=1'b0; c=1'b0; d=1'b0; #20;
	a=1'b1; b=1'b0; c=1'b0; d=1'b1; #20;
	a=1'b1; b=1'b0; c=1'b1; d=1'b0; #20;
	a=1'b1; b=1'b0; c=1'b1; d=1'b1; #20;
	a=1'b1; b=1'b1; c=1'b0; d=1'b0; #20;
	a=1'b1; b=1'b1; c=1'b0; d=1'b1; #20;
	a=1'b1; b=1'b1; c=1'b1; d=1'b0; #20;
	a=1'b1; b=1'b1; c=1'b1; d=1'b1; #20;
	$display ("TEST SUCESSFULL");
end
endmodule
